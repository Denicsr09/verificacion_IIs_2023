package my_package;
  parameter pckg_sz = 40;
  parameter fifo_depth = 11;
  parameter num_transacciones = 6;
endpackage
