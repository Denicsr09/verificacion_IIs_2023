`define ROWS 4
`define COLUMS 4
`define pckg_sz 40
`define deep_fifo 4
`define num_transaciones 3
