`define pckg_sz 49
`define deep_fifo 3
`define num_transaciones  668
`define ROWS 4
`define COLUMS 4
