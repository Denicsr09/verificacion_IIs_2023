package my_package;
  parameter pckg_sz = 45;
  parameter fifo_depth = 7;
  parameter num_transacciones = 10;
endpackage
