`define pckg_size 46
`define deep_fifo 5
`define num_transacciones 729
`define ROWS 4
`define COLUMS 4
