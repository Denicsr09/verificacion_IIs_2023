`define ROWS 4
`define COLUMS 4
`define pckg_sz 40

